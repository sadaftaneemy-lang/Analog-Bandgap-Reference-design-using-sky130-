*general purpose bandgap reference circuit avsdbgp_3v3- technology: sky130

.options savecurrents

* Load Sky130 device models
.lib "/home/sadaf/Desktop/Majorproject2025/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/models/sky130.lib.spice" tt
*.include "/home/sadaf/Desktop/Majorproject2025/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/models/sky130.lib.spice"
*BGR circuit

XM1 A C VDD VDD sky130_fd_pr__pfet_g5v0d10v5 l=5 w=20
XM2 C C VDD VDD sky130_fd_pr__pfet_g5v0d10v5 l=5 w=20
XM3 H C VDD VDD sky130_fd_pr__pfet_g5v0d10v5 l=5 w=20
XM4 A A B GND sky130_fd_pr__nfet_g5v0d10v5 l=5 w=20
XM5 C A D GND sky130_fd_pr__nfet_g5v0d10v5 l=5 w=20

X6 GND GND I GND sky130_fd_pr__pnp_05v5_W3p40L3p40 M=1
X7 GND GND E GND sky130_fd_pr__pnp_05v5_W3p40L3p40 M=8
X8 GND GND F GND sky130_fd_pr__pnp_05v5_W3p40L3p40 M=1

*Start-up  circuit

XM9 C G GND GND sky130_fd_pr__nfet_g5v0d10v5 l=5 w=20
XM10 G A GND GND sky130_fd_pr__nfet_g5v0d10v5 l=1 w=20

*Enable circuit

XM11 B En Vx GND sky130_fd_pr__nfet_g5v0d10v5 l=5 w=20
XM12 D En Vy GND sky130_fd_pr__nfet_g5v0d10v5 l=5 w=20
XM13 H En Vz GND sky130_fd_pr__nfet_g5v0d10v5 l=5 w=20
XM14 K En G GND sky130_fd_pr__nfet_g5v0d10v5 l=5 w=20

R1 J E 2K
R2 F Vref 2K
R3 VDDA Vw 2K
RL GND Vref 100MEG

V1 Vw K DC 0V
V2 Vx I DC 0V
V3 Vy J DC 0V
V4 Vz Vref DC 0V

VDDA VDD GND DC 3.3V
VD En GND DC 3.3V

.dc temp -40 140 0.

.control
run
plot v(Vref) v(f) v(Vref,f)
plot v(Vref)
plot v(f)
.endc

.end




